module dictionary

interface Dictionary {
	lookup(string) ?Result
}
