module anki

pub struct Card {
pub:
	front string
	back  string
}
